module AND (
    input wire a,
    input wire b,
    output reg y
);

    assign y = a & b;
    
endmodule

